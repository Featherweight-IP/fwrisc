
`include "fwrisc_formal_opcode_defines.svh"

`itype_xor(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`rtype_xor(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`rtype_sll(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`rtype_slt(idata, $anyconst, $anyconst, $anyconst);
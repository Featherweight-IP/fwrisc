


module fwrisc_decode_formal_checker(
		// TODO: fill in port list
		);
	
endmodule
		
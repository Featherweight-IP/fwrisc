
`include "fwrisc_formal_opcode_defines.svh"

`rtype_add(idata, $anyconst, $anyconst, $anyconst);
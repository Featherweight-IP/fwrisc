
`include "fwrisc_formal_opcode_defines.svh"

`rtype_sra(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`itype_sltu(idata, $anyconst, $anyconst, $anyconst);
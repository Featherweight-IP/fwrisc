
`include "fwrisc_formal_opcode_defines.svh"

`jalr(idata, $anyconst, $anyconst, $anyconst);
// `jal(idata, 4, $anyconst);
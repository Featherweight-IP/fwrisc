/****************************************************************************
 * rv32_tracer_bfm.sv
 ****************************************************************************/

/**
 * Module: rv32_tracer_bfm
 * 
 * TODO: Add interface documentation
 */
module rv32_tracer_bfm(
		input				clock,
		input				reset,
		input [31:0]		pc,
		input [31:0]		insn,
		input [31:0]		rs1,
		input [31:0]		rs2,
		input [31:0]		rt
		);

	

endmodule




`include "fwrisc_formal_opcode_defines.svh"

`utype_lui(idata, $anyconst, $anyconst);
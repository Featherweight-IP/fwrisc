
`include "fwrisc_formal_opcode_defines.svh"

`rtype_sub(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`jal(idata, $anyconst, $anyconst);


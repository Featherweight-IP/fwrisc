
`include "fwrisc_formal_opcode_defines.svh"

`rtype_or(idata, $anyconst, $anyconst, $anyconst);



module fwrisc_mem_checker(
		// TODO: fill in port list
		);
	
endmodule
		
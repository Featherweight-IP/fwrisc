
`include "fwrisc_formal_opcode_defines.svh"

`rtype_and(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`itype_add(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`itype_sll(idata, $anyconst, $anyconst, $anyconst);
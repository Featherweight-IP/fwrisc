
`include "fwrisc_formal_opcode_defines.svh"

`rtype_sltu(idata, $anyconst, $anyconst, $anyconst);
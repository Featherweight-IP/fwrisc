
`include "fwrisc_formal_opcode_defines.svh"

`rtype_srl(idata, $anyconst, $anyconst, $anyconst);
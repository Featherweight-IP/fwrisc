
`include "fwrisc_formal_opcode_defines.svh"

`itype_or(idata, $anyconst, $anyconst, $anyconst);

`include "fwrisc_formal_opcode_defines.svh"

`itype_slt(idata, $anyconst, $anyconst, $anyconst);
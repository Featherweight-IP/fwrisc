


module fwrisc_fetch_formal_test(
		// TODO: specify portlist
		);
	

endmodule